module simplified_sha256_part2 #(
	parameter integer NUM_OF_WORDS = 16)
	
(input logic  clk, reset_n, start,
 output logic done,
 output logic [31:0] mem_write_data[8], // changed mem_write_data to a vector
 input logic [31:0] mem_read_data[16], // changed mem_read_data to a vector, meant to connect to sha256_in
 input logic [31:0] hash[8]); //h0 to h7 controlled by hash vector

// FSM state variables 
enum logic [2:0] {IDLE, READ, BLOCK, COMPUTE, WRITE} state;

// Local variables
logic [31:0] w[16];
logic [31:0] message[16];
logic [31:0] wt;
logic [31:0] h0, h1, h2, h3, h4, h5, h6, h7;
logic [31:0] a, b, c, d, e, f, g, h;
logic [ 7:0] i, j;
logic [ 7:0] num_blocks;
logic [7:0]  curr_block;
logic [15:0] cur_addr;
logic [31:0] cur_write_data[8];
logic [512:0] memory_block;

// SHA256 K constants
parameter int k[0:63] = '{
   32'h428a2f98,32'h71374491,32'hb5c0fbcf,32'he9b5dba5,32'h3956c25b,32'h59f111f1,32'h923f82a4,32'hab1c5ed5,
   32'hd807aa98,32'h12835b01,32'h243185be,32'h550c7dc3,32'h72be5d74,32'h80deb1fe,32'h9bdc06a7,32'hc19bf174,
   32'he49b69c1,32'hefbe4786,32'h0fc19dc6,32'h240ca1cc,32'h2de92c6f,32'h4a7484aa,32'h5cb0a9dc,32'h76f988da,
   32'h983e5152,32'ha831c66d,32'hb00327c8,32'hbf597fc7,32'hc6e00bf3,32'hd5a79147,32'h06ca6351,32'h14292967,
   32'h27b70a85,32'h2e1b2138,32'h4d2c6dfc,32'h53380d13,32'h650a7354,32'h766a0abb,32'h81c2c92e,32'h92722c85,
   32'ha2bfe8a1,32'ha81a664b,32'hc24b8b70,32'hc76c51a3,32'hd192e819,32'hd6990624,32'hf40e3585,32'h106aa070,
   32'h19a4c116,32'h1e376c08,32'h2748774c,32'h34b0bcb5,32'h391c0cb3,32'h4ed8aa4a,32'h5b9cca4f,32'h682e6ff3,
   32'h748f82ee,32'h78a5636f,32'h84c87814,32'h8cc70208,32'h90befffa,32'ha4506ceb,32'hbef9a3f7,32'hc67178f2
};


assign num_blocks = 1; // should only support one block
assign wt = w[0];
assign mem_write_data = cur_write_data;

function logic [15:0] determine_num_blocks(input logic [31:0] size);

  determine_num_blocks = size / 512 + (size % 512 != 0);

endfunction


// SHA256 hash round
function logic [255:0] sha256_op(input logic [31:0] a, b, c, d, e, f, g, h, w,
                                 input logic [7:0] t);
    logic [31:0] S1, S0, ch, maj, t1, t2; // internal signals
begin
    S1 = rightrotate(e, 6) ^ rightrotate(e, 11) ^ rightrotate(e, 25);
    ch = (e & f) ^ (~e & g);
    t1 = h + S1 + ch + k[t] + w;
    S0 = rightrotate(a,2) ^ rightrotate(a,13) ^ rightrotate(a,22);
    maj = (a & b) ^ (a & c) ^ (b & c);
    t2 = S0 + maj;
    sha256_op = {t1 + t2, a, b, c, d + t1, e, f, g};
end
endfunction

function logic [31:0] rightrotate(input logic [31:0] x,
                                  input logic [ 7:0] r);
   rightrotate = (x >> r) | (x << (32 - r));
endfunction

function logic [31:0] wtnew;
	logic[31:0] s0,s1;
	begin
		s0 = rightrotate(w[1],7)^rightrotate(w[1],18)^(w[1]>>3);
		s1 = rightrotate(w[14],17)^rightrotate(w[14],19)^(w[14]>>10);
		wtnew = w[0] + s0 + w[9] + s1;
	end
endfunction

always_ff @(posedge clk, negedge reset_n)
begin
  if (!reset_n) begin
    state <= IDLE;
  end 
  else case (state)
    // Initialize hash values h0 to h7 and a to h, other variables and memory we, address offset, etc
    IDLE: begin 
       if(start) begin
			h0 <= hash[0]; // starting h seed based on hash vector, so we can modify it from outside
			h1 <= hash[1];
			h2 <= hash[2];
			h3 <= hash[3];
			h4 <= hash[4];
			h5 <= hash[5];
			h6 <= hash[6];
			h7 <= hash[7];
			curr_block <= 0;
			state <= READ;
       end else begin
			state <= IDLE;
		 end
    end
	 
	 READ: begin
		for (int n = 0; n < 16; n++)
		  message[n] <= mem_read_data[n];
		state <= BLOCK;
     end

    BLOCK: begin
			if (curr_block == num_blocks) begin
				state <= WRITE;
			end else begin
				for (int l = 0; l < 16; l++) begin
					w[l] <= message[l];
				end
				a = h0;
				b = h1;
				c = h2;
				d = h3;
				e = h4;
				f = h5;
				g = h6;
				h = h7;
				i <= 0;
				state <= COMPUTE;
			end
    end

    COMPUTE: begin
        if (i < 64) begin
			for (int m = 0; m < 15; m++) begin
				w[m] <= w[m+1];
			end
			w[15] <= wtnew;
			{a,b,c,d,e,f,g,h} <= sha256_op(a,b,c,d,e,f,g,h,wt,i);
			i <= i + 1;
			state <= COMPUTE;
        end else begin
			h0 <= h0 + a;
			h1 <= h1 + b;
			h2 <= h2 + c;
			h3 <= h3 + d;
			h4 <= h4 + e;
			h5 <= h5 + f;
			h6 <= h6 + g;
			h7 <= h7 + h;
			curr_block <= curr_block + 1;
         state <= BLOCK;
		  end
    end

    WRITE: begin
			cur_write_data[0] <= h0;
			cur_write_data[1] <= h1;
			cur_write_data[2] <= h2;            
			cur_write_data[3] <= h3;             
			cur_write_data[4] <= h4;             
			cur_write_data[5] <= h5;             
			cur_write_data[6] <= h6;          
			cur_write_data[7] <= h7;
			state <= IDLE;
    end
	 
	 endcase
  end
  
assign done = (state == IDLE);

endmodule
